module simple_memory#(
	parameter [ 31:0] pWords = 32'd128
)(
	input wire iwClk,
	input wire iwnRst,

	input wire [31:0]iwReadAddr,
	input wire [31:0]iwWriteAddr,
	input wire [31:0]iwWriteData,
	input wire [3:0]iwWstrb,

	output wire [31:0]owReadData,
	output wire [31:0]owLastData
);
reg [7:0]rMemory[0:pWords * 4 - 1];

assign owReadData[7:0] = rMemory[iwReadAddr];
assign owReadData[15:8] = rMemory[iwReadAddr + 1];
assign owReadData[23:16] = rMemory[iwReadAddr + 2];
assign owReadData[31:24] = rMemory[iwReadAddr + 3];

assign owLastData[7:0] = rMemory[pWords * 4 - 4];
assign owLastData[15:8] = rMemory[pWords * 4 - 3];
assign owLastData[23:16] = rMemory[pWords * 4 - 2];
assign owLastData[31:24] = rMemory[pWords * 4 - 1];

initial begin
	`include "simple_memory_rom.v"
end

always @(posedge iwClk or negedge iwnRst) begin
	if (!iwnRst) begin
		rMemory[pWords * 4 - 1] = 0;
		rMemory[pWords * 4 - 2] = 0;
		rMemory[pWords * 4 - 3] = 0;
		rMemory[pWords * 4 - 4] = 0;
	end else begin
		if (iwWstrb & 4'b1)
			rMemory[iwWriteAddr] = iwWriteData[7:0];
		if (iwWstrb & 4'b10)
			rMemory[iwWriteAddr + 1] = iwWriteData[15:8];
		if (iwWstrb & 4'b10)
			rMemory[iwWriteAddr + 2] = iwWriteData[23:16];
		if (iwWstrb & 4'b1000)
			rMemory[iwWriteAddr + 3] = iwWriteData[31:24];
	end
end

endmodule
